module inverter(input a, output b);
        assign b = ~a;
endmodule
